// (c) Copyright 2007 Actel Corporation
// Rev:                 2.1 15Mar107 AS - Production
module
CORESPI
#
(
parameter
FAMILY
=
17
,
parameter
USE_MASTER
=
1
,
parameter
USE_SLAVE
=
1
)
(
input
PCLK,
input
PRESETN,
output
m_sck,
input
m_miso,
output
m_mosi,
output
[
7
:
0
]
m_ss,
input
s_sck,
output
s_miso,
input
s_mosi,
input
s_ss,
output
enable_master,
output
enable_slave,
output
interrupt,
output
tx_reg_empty,
output
rx_data_ready,
input
PSEL,
input
PENABLE,
input
PWRITE,
input
[
3
:
0
]
PADDR,
input
[
7
:
0
]
PWDATA,
output
[
7
:
0
]
PRDATA
)
;
wire
[
7
:
0
]
CSPIO
;
wire
[
7
:
0
]
CSPII
;
wire
[
1
:
0
]
CSPIl
;
wire
CSPIOI
;
wire
CSPIII
;
assign
CSPIOI
=
(
PWRITE
&&
PSEL
&&
PENABLE
)
;
assign
CSPIII
=
(
~
PWRITE
&&
PSEL
&&
PENABLE
)
;
assign
CSPIO
=
PWDATA
;
assign
PRDATA
=
CSPII
;
assign
CSPIl
=
PADDR
[
3
:
2
]
;
CSPIlI
#
(
.USE_MASTER
(
USE_MASTER
)
,
.USE_SLAVE
(
USE_SLAVE
)
)
CSPIOl
(
.sysclk
(
PCLK
)
,
.nreset
(
PRESETN
)
,
.m_sck
(
m_sck
)
,
.m_miso
(
m_miso
)
,
.m_mosi
(
m_mosi
)
,
.m_ss
(
m_ss
)
,
.s_sck
(
s_sck
)
,
.s_miso
(
s_miso
)
,
.s_mosi
(
s_mosi
)
,
.s_ss
(
s_ss
)
,
.enable_master
(
enable_master
)
,
.enable_slave
(
enable_slave
)
,
.CSPIIl
(
CSPIO
)
,
.CSPIll
(
CSPII
)
,
.CSPIO0
(
CSPIl
)
,
.CSPII0
(
CSPIOI
)
,
.CSPIl0
(
CSPIII
)
,
.interrupt
(
interrupt
)
,
.tx_reg_empty
(
tx_reg_empty
)
,
.rx_data_ready
(
rx_data_ready
)
)
;
endmodule
