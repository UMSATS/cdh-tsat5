// (c) Copyright 2005 Actel Corporation
// Rev:                 2.1 24Jan05 TFB - Production
`timescale 1ns/1ps
module
spi_master
(
sysclk
,
nreset
,
enable
,
sck
,
miso
,
mosi
,
ss
,
cpol
,
cpha
,
clocksel
,
rx_data_reg
,
rx_data_ready
,
rx_reg_re
,
tx_data_reg
,
tx_reg_empty
,
busy
,
tx_reg_we
,
clear_error
,
rx_error
)
;
input
sysclk
;
input
nreset
;
input
enable
;
output
sck
;
input
miso
;
output
mosi
;
output
ss
;
input
cpol
;
input
cpha
;
input
[
2
:
0
]
clocksel
;
output
[
7
:
0
]
rx_data_reg
;
output
rx_data_ready
;
input
rx_reg_re
;
input
[
7
:
0
]
tx_data_reg
;
output
tx_reg_empty
;
output
busy
;
input
tx_reg_we
;
input
clear_error
;
output
rx_error
;
wire
sck
;
wire
ss
;
wire
rx_data_ready
;
wire
tx_reg_empty
;
wire
busy
;
wire
rx_error
;
reg
mosi
;
reg
[
7
:
0
]
rx_data_reg
;
parameter
[
3
:
0
]
CSPIOO0
=
0
,
CSPIIO0
=
1
,
CSPIlO0
=
2
,
CSPIOI0
=
3
,
CSPIII0
=
4
,
D3
=
5
,
D2
=
6
,
D1
=
7
,
D0
=
8
,
CSPIlI0
=
9
,
CSPIOl0
=
10
;
reg
[
3
:
0
]
CSPIIl0
;
reg
[
3
:
0
]
CSPIll0
;
reg
CSPIO00
;
reg
CSPII00
;
wire
CSPIl00
;
reg
CSPIO10
;
reg
CSPII10
;
reg
CSPIl10
;
reg
CSPIlOl
;
reg
[
7
:
0
]
CSPIOO1
;
reg
CSPIIO1
;
reg
CSPIlO1
;
reg
[
7
:
0
]
CSPIOI1
;
reg
[
7
:
0
]
CSPIII1
;
reg
CSPIlI1
;
reg
CSPIOl1
;
reg
CSPIIl1
;
reg
CSPIll1
;
reg
CSPIO01
;
reg
CSPII01
;
reg
CSPIl01
;
reg
CSPIO11
;
reg
CSPII11
;
wire
CSPIl11
;
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIOO1
<=
{
8
{
1
'b
0
}
}
;
CSPIO00
<=
1
'b
0
;
CSPII00
<=
1
'b
0
;
end
else
begin
if
(
enable
==
1
'b
1
)
begin
CSPIOO1
<=
CSPIOO1
+
8
'b
00000001
;
end
case
(
clocksel
)
3
'b
000
:
begin
CSPIO00
<=
CSPIOO1
[
0
]
;
end
3
'b
001
:
begin
CSPIO00
<=
CSPIOO1
[
1
]
;
end
3
'b
010
:
begin
CSPIO00
<=
CSPIOO1
[
2
]
;
end
3
'b
011
:
begin
CSPIO00
<=
CSPIOO1
[
3
]
;
end
3
'b
100
:
begin
CSPIO00
<=
CSPIOO1
[
4
]
;
end
3
'b
101
:
begin
CSPIO00
<=
CSPIOO1
[
5
]
;
end
3
'b
110
:
begin
CSPIO00
<=
CSPIOO1
[
6
]
;
end
3
'b
111
:
begin
CSPIO00
<=
CSPIOO1
[
7
]
;
end
default
:
begin
CSPIO00
<=
CSPIOO1
[
0
]
;
end
endcase
CSPII00
<=
CSPIO00
;
end
end
assign
CSPIl00
=
(
cpha
==
1
'b
1
&
cpol
==
1
'b
0
)
?
CSPIll1
&
CSPII00
:
(
cpha
==
1
'b
1
&
cpol
==
1
'b
1
)
?
~
(
CSPIll1
&
CSPII00
)
:
(
cpha
==
1
'b
0
&
cpol
==
1
'b
0
)
?
CSPIll1
&
(
~
CSPII00
)
:
~
(
CSPIll1
&
(
~
CSPII00
)
)
;
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIO10
<=
1
'b
0
;
end
else
begin
CSPIO10
<=
CSPIl00
;
end
end
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIl10
<=
1
'b
1
;
end
else
begin
CSPIl10
<=
CSPII10
;
end
end
assign
sck
=
CSPIO10
;
assign
ss
=
CSPIl10
;
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIIl0
<=
CSPIOO0
;
end
else
begin
if
(
enable
==
1
'b
1
)
begin
CSPIIl0
<=
CSPIll0
;
end
else
begin
CSPIIl0
<=
CSPIOO0
;
end
end
end
always
@
(
CSPIIl0
or
CSPIIO1
or
CSPIO00
or
CSPII00
)
begin
CSPIlO1
<=
1
'b
0
;
CSPIlI1
<=
1
'b
0
;
CSPIOl1
<=
1
'b
0
;
CSPII10
<=
1
'b
1
;
CSPIll1
<=
1
'b
0
;
CSPIO01
<=
1
'b
0
;
case
(
CSPIIl0
)
CSPIOO0
:
begin
if
(
CSPIIO1
==
1
'b
1
&
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
)
begin
CSPIlO1
<=
1
'b
1
;
CSPIll0
<=
CSPIOl0
;
end
else
begin
CSPIll0
<=
CSPIOO0
;
end
end
CSPIOl0
:
begin
CSPIOl1
<=
1
'b
1
;
if
(
CSPII00
==
1
'b
0
)
begin
CSPII10
<=
1
'b
0
;
if
(
CSPIO00
==
1
'b
1
)
begin
CSPIll0
<=
CSPIIO0
;
end
else
begin
CSPIll0
<=
CSPIOl0
;
end
end
else
begin
CSPIll0
<=
CSPIOl0
;
end
end
CSPIIO0
:
begin
CSPII10
<=
1
'b
0
;
CSPIll1
<=
1
'b
1
;
if
(
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
)
begin
CSPIlI1
<=
1
'b
1
;
CSPIll0
<=
CSPIlO0
;
end
else
begin
CSPIll0
<=
CSPIIO0
;
end
end
CSPIlO0
:
begin
CSPII10
<=
1
'b
0
;
CSPIll1
<=
1
'b
1
;
if
(
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
)
begin
CSPIlI1
<=
1
'b
1
;
CSPIll0
<=
CSPIOI0
;
end
else
begin
CSPIll0
<=
CSPIlO0
;
end
end
CSPIOI0
:
begin
CSPII10
<=
1
'b
0
;
CSPIll1
<=
1
'b
1
;
if
(
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
)
begin
CSPIlI1
<=
1
'b
1
;
CSPIll0
<=
CSPIII0
;
end
else
begin
CSPIll0
<=
CSPIOI0
;
end
end
CSPIII0
:
begin
CSPII10
<=
1
'b
0
;
CSPIll1
<=
1
'b
1
;
if
(
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
)
begin
CSPIlI1
<=
1
'b
1
;
CSPIll0
<=
D3
;
end
else
begin
CSPIll0
<=
CSPIII0
;
end
end
D3
:
begin
CSPII10
<=
1
'b
0
;
CSPIll1
<=
1
'b
1
;
if
(
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
)
begin
CSPIlI1
<=
1
'b
1
;
CSPIll0
<=
D2
;
end
else
begin
CSPIll0
<=
D3
;
end
end
D2
:
begin
CSPII10
<=
1
'b
0
;
CSPIll1
<=
1
'b
1
;
if
(
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
)
begin
CSPIlI1
<=
1
'b
1
;
CSPIll0
<=
D1
;
end
else
begin
CSPIll0
<=
D2
;
end
end
D1
:
begin
CSPII10
<=
1
'b
0
;
CSPIll1
<=
1
'b
1
;
if
(
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
)
begin
CSPIlI1
<=
1
'b
1
;
CSPIll0
<=
D0
;
end
else
begin
CSPIll0
<=
D1
;
end
end
D0
:
begin
CSPII10
<=
1
'b
0
;
CSPIll1
<=
1
'b
1
;
if
(
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
)
begin
CSPIlI1
<=
1
'b
1
;
CSPIll0
<=
CSPIlI0
;
end
else
begin
CSPIll0
<=
D0
;
end
end
CSPIlI0
:
begin
if
(
CSPII00
==
1
'b
1
)
begin
CSPII10
<=
1
'b
0
;
CSPIll0
<=
CSPIlI0
;
end
else
begin
CSPIO01
<=
1
'b
1
;
CSPII10
<=
1
'b
1
;
if
(
CSPIIO1
==
1
'b
1
&
CSPIO00
==
1
'b
1
)
begin
CSPIlO1
<=
1
'b
1
;
CSPIll0
<=
CSPIOl0
;
end
else
begin
CSPIll0
<=
CSPIOO0
;
end
end
end
endcase
end
always
@
(
CSPII10
or
CSPIl00
or
CSPIO10
or
cpol
or
cpha
)
begin
if
(
CSPII10
==
1
'b
0
)
begin
if
(
(
cpol
^
cpha
)
==
1
'b
0
)
begin
CSPIO11
<=
CSPIl00
&
(
~
CSPIO10
)
;
end
else
begin
CSPIO11
<=
(
~
CSPIl00
)
&
CSPIO10
;
end
end
else
begin
CSPIO11
<=
1
'b
0
;
end
end
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPII11
<=
1
'b
0
;
end
else
begin
CSPII11
<=
CSPIO11
;
end
end
assign
CSPIl11
=
(
clocksel
==
3
'b
000
)
?
CSPII11
:
CSPIO11
;
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIII1
<=
{
8
{
1
'b
0
}
}
;
end
else
begin
if
(
CSPIl11
==
1
'b
1
)
begin
CSPIII1
[
0
]
<=
miso
;
CSPIII1
[
7
:
1
]
<=
CSPIII1
[
6
:
0
]
;
end
end
end
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIOI1
<=
{
8
{
1
'b
0
}
}
;
mosi
<=
1
'b
0
;
end
else
begin
if
(
CSPIOl1
==
1
'b
1
)
begin
CSPIOI1
<=
tx_data_reg
;
end
else
if
(
CSPIlI1
==
1
'b
1
)
begin
CSPIOI1
[
7
:
1
]
<=
CSPIOI1
[
6
:
0
]
;
end
mosi
<=
CSPIOI1
[
7
]
;
end
end
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
rx_data_reg
<=
{
8
{
1
'b
0
}
}
;
end
else
begin
if
(
enable
==
1
'b
1
)
begin
if
(
CSPIO01
==
1
'b
1
)
begin
rx_data_reg
<=
CSPIII1
;
end
end
end
end
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIl01
<=
1
'b
0
;
CSPII01
<=
1
'b
0
;
end
else
begin
if
(
rx_reg_re
==
1
'b
1
)
begin
CSPIl01
<=
1
'b
0
;
end
else
if
(
clear_error
==
1
'b
1
)
begin
CSPII01
<=
1
'b
0
;
end
else
if
(
CSPIO01
==
1
'b
1
)
begin
if
(
CSPIl01
==
1
'b
1
)
begin
CSPII01
<=
1
'b
1
;
end
else
begin
CSPIl01
<=
1
'b
1
;
end
end
end
end
assign
rx_error
=
CSPII01
;
assign
rx_data_ready
=
CSPIl01
;
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIIO1
<=
1
'b
0
;
CSPIlOl
<=
1
'b
1
;
CSPIIl1
<=
1
'b
0
;
end
else
begin
if
(
tx_reg_we
==
1
'b
1
)
begin
CSPIIO1
<=
1
'b
1
;
CSPIlOl
<=
1
'b
0
;
end
else
if
(
CSPIlO1
==
1
'b
1
)
begin
CSPIIO1
<=
1
'b
0
;
end
else
if
(
CSPIOl1
==
1
'b
0
&
CSPIIl1
==
1
'b
1
)
begin
CSPIlOl
<=
1
'b
1
;
end
CSPIIl1
<=
CSPIOl1
;
end
end
assign
tx_reg_empty
=
CSPIlOl
;
assign
busy
=
(
CSPIl10
==
1
'b
0
|
(
~
CSPIlOl
)
==
1
'b
1
|
CSPIIl0
!=
CSPIOO0
)
?
1
'b
1
:
1
'b
0
;
endmodule
