// Copyright (c) 2009 Actel Corporation.  All rights reserved.
// Revision: CoreI2C v6.0  18Aug2009
// SVN Revision Information:
// SVN $Revision: 15634 $
`timescale 1ns/1ns
module
COREI2C
#
(
parameter
FAMILY
=
17
,
parameter
OPERATING_MODE
=
0
,
parameter
BAUD_RATE_FIXED
=
0
,
parameter
BAUD_RATE_VALUE
=
3
'b
000
,
parameter
BCLK_ENABLED
=
1
,
parameter
GLITCHREG_NUM
=
3
,
parameter
SMB_EN
=
0
,
parameter
IPMI_EN
=
1
,
parameter
FREQUENCY
=
30
,
parameter
FIXED_SLAVE0_ADDR_EN
=
0
,
parameter
FIXED_SLAVE0_ADDR_VALUE
=
8
'h
00
,
parameter
ADD_SLAVE1_ADDRESS_EN
=
1
,
parameter
FIXED_SLAVE1_ADDR_EN
=
0
,
parameter
FIXED_SLAVE1_ADDR_VALUE
=
8
'h
00
,
parameter
I2C_NUM
=
1
)
(
input
PRESETN,
input
PCLK,
input
BCLK,
input
PSEL,
input
PENABLE,
input
PWRITE,
input
[
8
:
0
]
PADDR,
input
[
7
:
0
]
PWDATA,
output
reg
[
7
:
0
]
PRDATA,
output
[
I2C_NUM
-
1
:
0
]
INT,
input
[
I2C_NUM
-
1
:
0
]
SCLI,
input
[
I2C_NUM
-
1
:
0
]
SDAI,
output
[
I2C_NUM
-
1
:
0
]
SCLO,
output
[
I2C_NUM
-
1
:
0
]
SDAO,
input
[
I2C_NUM
-
1
:
0
]
SMBALERT_NI,
output
[
I2C_NUM
-
1
:
0
]
SMBALERT_NO,
output
[
I2C_NUM
-
1
:
0
]
SMBA_INT,
input
[
I2C_NUM
-
1
:
0
]
SMBSUS_NI,
output
[
I2C_NUM
-
1
:
0
]
SMBSUS_NO,
output
[
I2C_NUM
-
1
:
0
]
SMBS_INT
)
;
function
[
31
:
0
]
CI2CO
;
input
integer
CI2CI
;
integer
CI2Cl
,
CI2COI
;
begin
CI2Cl
=
1
;
CI2COI
=
0
;
while
(
CI2Cl
<
CI2CI
)
begin
CI2Cl
=
CI2Cl
*
2
;
CI2COI
=
CI2COI
+
1
;
end
CI2CO
=
CI2COI
;
end
endfunction
parameter
[
4
:
0
]
CI2CII
=
5
'b
01100
;
parameter
[
7
:
0
]
CI2ClI
=
8
'b
00000000
;
parameter
[
4
:
0
]
CI2COl
=
5
'b
11100
;
parameter
[
7
:
0
]
CI2CIl
=
8
'b
00000000
;
wire
[
0
:
I2C_NUM
-
1
]
PSELi
;
wire
[
CI2CO
(
FREQUENCY
*
215
)
-
1
:
0
]
CI2Cll
=
(
FREQUENCY
*
215
)
;
reg
[
CI2CO
(
FREQUENCY
*
215
)
-
1
:
0
]
CI2CO0
;
wire
pulse_215us
;
reg
CI2CI0
;
reg
CI2Cl0
;
wire
BCLKe
;
reg
[
7
:
0
]
CI2CO1
;
wire
[
7
:
0
]
seradr0
;
reg
[
7
:
0
]
CI2CI1
;
wire
[
7
:
0
]
seradr1
;
wire
seradr1apb0
;
wire
[
7
:
0
]
CI2Cl1
[
0
:
I2C_NUM
-
1
]
;
assign
seradr1apb0
=
(
ADD_SLAVE1_ADDRESS_EN
==
1
)
?
CI2CI1
[
0
]
:
1
'b
0
;
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
begin
:
CI2COOI
if
(
PRESETN
==
1
'b
0
)
begin
CI2CO0
<=
0
;
end
else
begin
if
(
CI2CO0
==
0
)
begin
CI2CO0
<=
CI2Cll
;
end
else
begin
CI2CO0
<=
CI2CO0
-
1
;
end
end
end
assign
pulse_215us
=
(
(
CI2CO0
==
0
)
&&
(
(
IPMI_EN
==
1
)
||
(
SMB_EN
==
1
)
)
)
?
1
'b
1
:
1
'b
0
;
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
begin
:
CI2CIOI
if
(
PRESETN
==
1
'b
0
)
begin
CI2CI0
<=
1
'b
1
;
CI2Cl0
<=
1
'b
1
;
end
else
begin
CI2CI0
<=
BCLK
;
CI2Cl0
<=
CI2CI0
;
end
end
assign
BCLKe
=
BCLK_ENABLED
==
1
?
CI2CI0
&
~
CI2Cl0
:
1
'b
0
;
generate
begin
:
CI2ClOI
if
(
FIXED_SLAVE0_ADDR_EN
==
0
)
begin
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
begin
:
CI2COII
if
(
PRESETN
==
1
'b
0
)
begin
CI2CO1
<=
CI2ClI
;
end
else
begin
if
(
(
PENABLE
&&
PWRITE
&&
PSEL
)
&&
(
PADDR
[
4
:
0
]
==
CI2CII
)
)
begin
CI2CO1
<=
PWDATA
;
end
end
end
assign
seradr0
=
CI2CO1
;
end
else
begin
assign
seradr0
=
{
FIXED_SLAVE0_ADDR_VALUE
[
6
:
0
]
,
1
'b
0
}
;
end
end
endgenerate
generate
begin
:
CI2CIII
if
(
(
FIXED_SLAVE1_ADDR_EN
==
0
)
&&
(
ADD_SLAVE1_ADDRESS_EN
==
1
)
)
begin
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
begin
:
CI2ClII
if
(
PRESETN
==
1
'b
0
)
begin
CI2CI1
<=
CI2CIl
;
end
else
begin
if
(
(
PENABLE
&&
PWRITE
&&
PSEL
)
&&
(
PADDR
[
4
:
0
]
==
CI2COl
)
)
begin
CI2CI1
<=
PWDATA
;
end
end
end
assign
seradr1
=
CI2CI1
;
end
else
if
(
(
FIXED_SLAVE1_ADDR_EN
==
1
)
&&
(
ADD_SLAVE1_ADDRESS_EN
==
1
)
)
begin
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
begin
:
CI2ClII
if
(
PRESETN
==
1
'b
0
)
begin
CI2CI1
<=
{
7
'b
0
,
CI2CIl
[
0
]
}
;
end
else
begin
if
(
(
PENABLE
&&
PWRITE
&&
PSEL
)
&&
(
PADDR
[
4
:
0
]
==
CI2COl
)
)
begin
CI2CI1
<=
{
7
'b
0
,
PWDATA
[
0
]
}
;
end
end
end
assign
seradr1
=
{
FIXED_SLAVE1_ADDR_VALUE
[
6
:
0
]
,
CI2CI1
[
0
]
}
;
end
else
begin
assign
seradr1
=
8
'b
0
;
end
end
endgenerate
genvar
CI2COlI
;
generate
for
(
CI2COlI
=
0
;
CI2COlI
<=
(
I2C_NUM
-
1
)
;
CI2COlI
=
CI2COlI
+
1
)
begin
:
CI2CIlI
COREI2CREAL
#
(
.FAMILY
(
FAMILY
)
,
.OPERATING_MODE
(
OPERATING_MODE
)
,
.BAUD_RATE_FIXED
(
BAUD_RATE_FIXED
)
,
.BAUD_RATE_VALUE
(
BAUD_RATE_VALUE
)
,
.BCLK_ENABLED
(
BCLK_ENABLED
)
,
.GLITCHREG_NUM
(
GLITCHREG_NUM
)
,
.SMB_EN
(
SMB_EN
)
,
.IPMI_EN
(
IPMI_EN
)
,
.FREQUENCY
(
FREQUENCY
)
,
.FIXED_SLAVE0_ADDR_EN
(
FIXED_SLAVE0_ADDR_EN
)
,
.FIXED_SLAVE0_ADDR_VALUE
(
FIXED_SLAVE0_ADDR_VALUE
)
,
.ADD_SLAVE1_ADDRESS_EN
(
ADD_SLAVE1_ADDRESS_EN
)
,
.FIXED_SLAVE1_ADDR_EN
(
FIXED_SLAVE1_ADDR_EN
)
,
.FIXED_SLAVE1_ADDR_VALUE
(
FIXED_SLAVE1_ADDR_VALUE
)
)
ui2c
(
.pulse_215us
(
pulse_215us
)
,
.seradr0
(
seradr0
)
,
.seradr1apb0
(
seradr1apb0
)
,
.seradr1
(
seradr1
)
,
.PCLK
(
PCLK
)
,
.PRESETN
(
PRESETN
)
,
.BCLKe
(
BCLKe
)
,
.SCLI
(
SCLI
[
CI2COlI
]
)
,
.SDAI
(
SDAI
[
CI2COlI
]
)
,
.SCLO
(
SCLO
[
CI2COlI
]
)
,
.SDAO
(
SDAO
[
CI2COlI
]
)
,
.INT
(
INT
[
CI2COlI
]
)
,
.PWDATA
(
PWDATA
)
,
.PRDATA
(
CI2Cl1
[
CI2COlI
]
)
,
.PADDR
(
PADDR
[
4
:
0
]
)
,
.PSEL
(
PSELi
[
CI2COlI
]
)
,
.PENABLE
(
PENABLE
)
,
.PWRITE
(
PWRITE
)
,
.SMBALERT_NI
(
SMBALERT_NI
[
CI2COlI
]
)
,
.SMBALERT_NO
(
SMBALERT_NO
[
CI2COlI
]
)
,
.SMBA_INT
(
SMBA_INT
[
CI2COlI
]
)
,
.SMBSUS_NI
(
SMBSUS_NI
[
CI2COlI
]
)
,
.SMBSUS_NO
(
SMBSUS_NO
[
CI2COlI
]
)
,
.SMBS_INT
(
SMBS_INT
[
CI2COlI
]
)
)
;
end
endgenerate
genvar
CI2CI
;
generate
for
(
CI2CI
=
0
;
CI2CI
<=
(
I2C_NUM
-
1
)
;
CI2CI
=
CI2CI
+
1
)
begin
:
CI2CllI
assign
PSELi
[
CI2CI
]
=
PSEL
&
(
PADDR
[
8
:
5
]
==
CI2CI
)
;
end
endgenerate
generate
if
(
I2C_NUM
==
1
)
begin
:
CI2CO0I
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
2
)
begin
:
CI2CI0I
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
3
)
begin
:
CI2Cl0I
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
4
)
begin
:
CI2CO1I
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
5
)
begin
:
CI2CI1I
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
6
)
begin
:
CI2Cl1I
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
7
)
begin
:
CI2COOl
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
4
'h
6
:
PRDATA
=
CI2Cl1
[
6
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
8
)
begin
:
CI2CIOl
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
4
'h
6
:
PRDATA
=
CI2Cl1
[
6
]
;
4
'h
7
:
PRDATA
=
CI2Cl1
[
7
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
9
)
begin
:
CI2ClOl
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
4
'h
6
:
PRDATA
=
CI2Cl1
[
6
]
;
4
'h
7
:
PRDATA
=
CI2Cl1
[
7
]
;
4
'h
8
:
PRDATA
=
CI2Cl1
[
8
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
10
)
begin
:
CI2COIl
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
4
'h
6
:
PRDATA
=
CI2Cl1
[
6
]
;
4
'h
7
:
PRDATA
=
CI2Cl1
[
7
]
;
4
'h
8
:
PRDATA
=
CI2Cl1
[
8
]
;
4
'h
9
:
PRDATA
=
CI2Cl1
[
9
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
11
)
begin
:
CI2CIIl
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
4
'h
6
:
PRDATA
=
CI2Cl1
[
6
]
;
4
'h
7
:
PRDATA
=
CI2Cl1
[
7
]
;
4
'h
8
:
PRDATA
=
CI2Cl1
[
8
]
;
4
'h
9
:
PRDATA
=
CI2Cl1
[
9
]
;
4
'h
a
:
PRDATA
=
CI2Cl1
[
10
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
12
)
begin
:
CI2ClIl
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
4
'h
6
:
PRDATA
=
CI2Cl1
[
6
]
;
4
'h
7
:
PRDATA
=
CI2Cl1
[
7
]
;
4
'h
8
:
PRDATA
=
CI2Cl1
[
8
]
;
4
'h
9
:
PRDATA
=
CI2Cl1
[
9
]
;
4
'h
a
:
PRDATA
=
CI2Cl1
[
10
]
;
4
'h
b
:
PRDATA
=
CI2Cl1
[
11
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
13
)
begin
:
CI2COll
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
4
'h
6
:
PRDATA
=
CI2Cl1
[
6
]
;
4
'h
7
:
PRDATA
=
CI2Cl1
[
7
]
;
4
'h
8
:
PRDATA
=
CI2Cl1
[
8
]
;
4
'h
9
:
PRDATA
=
CI2Cl1
[
9
]
;
4
'h
a
:
PRDATA
=
CI2Cl1
[
10
]
;
4
'h
b
:
PRDATA
=
CI2Cl1
[
11
]
;
4
'h
c
:
PRDATA
=
CI2Cl1
[
12
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
14
)
begin
:
CI2CIll
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
4
'h
6
:
PRDATA
=
CI2Cl1
[
6
]
;
4
'h
7
:
PRDATA
=
CI2Cl1
[
7
]
;
4
'h
8
:
PRDATA
=
CI2Cl1
[
8
]
;
4
'h
9
:
PRDATA
=
CI2Cl1
[
9
]
;
4
'h
a
:
PRDATA
=
CI2Cl1
[
10
]
;
4
'h
b
:
PRDATA
=
CI2Cl1
[
11
]
;
4
'h
c
:
PRDATA
=
CI2Cl1
[
12
]
;
4
'h
d
:
PRDATA
=
CI2Cl1
[
13
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
15
)
begin
:
CI2Clll
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
4
'h
6
:
PRDATA
=
CI2Cl1
[
6
]
;
4
'h
7
:
PRDATA
=
CI2Cl1
[
7
]
;
4
'h
8
:
PRDATA
=
CI2Cl1
[
8
]
;
4
'h
9
:
PRDATA
=
CI2Cl1
[
9
]
;
4
'h
a
:
PRDATA
=
CI2Cl1
[
10
]
;
4
'h
b
:
PRDATA
=
CI2Cl1
[
11
]
;
4
'h
c
:
PRDATA
=
CI2Cl1
[
12
]
;
4
'h
d
:
PRDATA
=
CI2Cl1
[
13
]
;
4
'h
e
:
PRDATA
=
CI2Cl1
[
14
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
generate
if
(
I2C_NUM
==
16
)
begin
:
CI2CO0l
always
@
*
begin
case
(
PADDR
[
8
:
5
]
)
4
'h
0
:
PRDATA
=
CI2Cl1
[
0
]
;
4
'h
1
:
PRDATA
=
CI2Cl1
[
1
]
;
4
'h
2
:
PRDATA
=
CI2Cl1
[
2
]
;
4
'h
3
:
PRDATA
=
CI2Cl1
[
3
]
;
4
'h
4
:
PRDATA
=
CI2Cl1
[
4
]
;
4
'h
5
:
PRDATA
=
CI2Cl1
[
5
]
;
4
'h
6
:
PRDATA
=
CI2Cl1
[
6
]
;
4
'h
7
:
PRDATA
=
CI2Cl1
[
7
]
;
4
'h
8
:
PRDATA
=
CI2Cl1
[
8
]
;
4
'h
9
:
PRDATA
=
CI2Cl1
[
9
]
;
4
'h
a
:
PRDATA
=
CI2Cl1
[
10
]
;
4
'h
b
:
PRDATA
=
CI2Cl1
[
11
]
;
4
'h
c
:
PRDATA
=
CI2Cl1
[
12
]
;
4
'h
d
:
PRDATA
=
CI2Cl1
[
13
]
;
4
'h
e
:
PRDATA
=
CI2Cl1
[
14
]
;
4
'h
f
:
PRDATA
=
CI2Cl1
[
15
]
;
default
:
PRDATA
=
8
'h
00
;
endcase
end
end
endgenerate
endmodule
