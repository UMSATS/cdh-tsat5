// (c) Copyright 2005 Actel Corporation
// Rev:                 2.1 24Jan05 TFB - Production
`timescale 1ns/1ps
module
spi_slave
(
sysclk
,
nreset
,
enable
,
sck
,
miso
,
mosi
,
ss
,
cpol
,
cpha
,
rx_data_reg
,
rx_data_ready
,
rx_reg_re
,
tx_data_reg
,
tx_reg_we
,
tx_reg_empty
,
clear_error
,
rx_error
)
;
input
sysclk
;
input
nreset
;
input
enable
;
input
sck
;
output
miso
;
input
mosi
;
input
ss
;
input
cpol
;
input
cpha
;
output
[
7
:
0
]
rx_data_reg
;
output
rx_data_ready
;
input
rx_reg_re
;
input
[
7
:
0
]
tx_data_reg
;
input
tx_reg_we
;
output
tx_reg_empty
;
input
clear_error
;
output
rx_error
;
wire
miso
;
wire
rx_data_ready
;
wire
rx_error
;
reg
[
7
:
0
]
rx_data_reg
;
reg
tx_reg_empty
;
reg
CSPIO00
;
reg
CSPII00
;
reg
CSPIOOOI
;
reg
CSPIIOOI
;
reg
CSPII10
;
reg
CSPIlOOI
;
reg
CSPIOIOI
;
reg
[
7
:
0
]
CSPIIIOI
;
wire
CSPIlIOI
;
reg
CSPIl01
;
reg
CSPII01
;
reg
[
3
:
0
]
CSPIOlOI
;
reg
CSPIIlOI
;
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIO00
<=
1
'b
0
;
CSPII00
<=
1
'b
0
;
CSPIOOOI
<=
1
'b
0
;
CSPIIOOI
<=
1
'b
0
;
CSPII10
<=
1
'b
1
;
CSPIlOOI
<=
1
'b
1
;
end
else
begin
if
(
enable
==
1
'b
1
)
begin
CSPIIOOI
<=
mosi
;
CSPIlOOI
<=
ss
;
if
(
cpol
==
1
'b
0
&
cpha
==
1
'b
0
)
begin
CSPIO00
<=
sck
;
end
else
if
(
cpol
==
1
'b
0
&
cpha
==
1
'b
1
)
begin
CSPIO00
<=
~
sck
;
end
else
if
(
cpol
==
1
'b
1
&
cpha
==
1
'b
0
)
begin
CSPIO00
<=
~
sck
;
end
else
begin
CSPIO00
<=
sck
;
end
CSPII00
<=
CSPIO00
;
CSPIOOOI
<=
CSPIIOOI
;
CSPII10
<=
CSPIlOOI
;
end
else
begin
CSPIlOOI
<=
1
'b
1
;
end
end
end
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIIIOI
<=
{
8
{
1
'b
0
}
}
;
CSPIIlOI
<=
1
'b
0
;
end
else
begin
if
(
CSPII10
==
1
'b
1
)
begin
CSPIIIOI
<=
tx_data_reg
;
end
else
if
(
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
)
begin
CSPIIIOI
[
0
]
<=
CSPIOOOI
;
CSPIIIOI
[
7
:
1
]
<=
CSPIIIOI
[
6
:
0
]
;
end
if
(
CSPIO00
==
1
'b
1
&
CSPII00
==
1
'b
0
&
CSPII10
==
1
'b
0
)
begin
CSPIIlOI
<=
1
'b
1
;
end
else
begin
CSPIIlOI
<=
1
'b
0
;
end
end
end
assign
miso
=
CSPIIIOI
[
7
]
;
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIOlOI
<=
4
'b
0000
;
end
else
begin
if
(
CSPII10
==
1
'b
1
|
CSPIOlOI
==
4
'b
1000
)
begin
CSPIOlOI
<=
4
'b
0000
;
end
else
if
(
CSPIIlOI
==
1
'b
1
)
begin
CSPIOlOI
<=
CSPIOlOI
+
4
'b
0001
;
end
end
end
assign
CSPIlIOI
=
CSPIOlOI
[
3
]
&
(
~
CSPIOlOI
[
2
]
)
&
(
~
CSPIOlOI
[
1
]
)
&
(
~
CSPIOlOI
[
0
]
)
;
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
tx_reg_empty
<=
1
'b
1
;
CSPIOIOI
<=
1
'b
0
;
end
else
begin
if
(
CSPII10
==
1
'b
0
&
CSPIOIOI
==
1
'b
1
)
begin
tx_reg_empty
<=
1
'b
1
;
end
else
if
(
tx_reg_we
==
1
'b
1
)
begin
tx_reg_empty
<=
1
'b
0
;
end
CSPIOIOI
<=
CSPII10
;
end
end
assign
rx_data_ready
=
CSPIl01
;
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
CSPIl01
<=
1
'b
0
;
CSPII01
<=
1
'b
0
;
end
else
begin
if
(
clear_error
==
1
'b
1
)
begin
CSPIl01
<=
1
'b
0
;
CSPII01
<=
1
'b
0
;
end
else
if
(
CSPIlIOI
==
1
'b
1
)
begin
if
(
CSPIl01
==
1
'b
1
)
begin
CSPII01
<=
1
'b
1
;
end
CSPIl01
<=
1
'b
1
;
end
else
if
(
rx_reg_re
==
1
'b
1
)
begin
CSPIl01
<=
1
'b
0
;
end
end
end
assign
rx_error
=
CSPII01
;
always
@
(
posedge
sysclk
or
negedge
nreset
)
begin
if
(
nreset
==
1
'b
0
)
begin
rx_data_reg
<=
8
'b
00000000
;
end
else
begin
if
(
enable
==
1
'b
1
)
begin
if
(
CSPIlIOI
==
1
'b
1
)
begin
rx_data_reg
<=
CSPIIIOI
;
end
end
end
end
endmodule
